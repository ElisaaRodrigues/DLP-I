---------------------
-- FILE my_pkg.vhd --
---------------------
library ieee;
use ieee.std_logic_1164.all;
 
package my_pkg is
	type a_slv	is array(natural range <>) of std_logic_vector (3 downto 0);
end package;